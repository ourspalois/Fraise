module MC_64x64_FULL_upd (
    input logic [63:0] CBL, 
    input logic [63:0] CBLEN, 
    input logic [63:0] CSL,
    input logic [63:0] DIN,
    input logic [63:0] DINb,
    
    input logic [31:0] CWLE,
    input logic [31:0] CWLO,

    input logic [63:0] DOUT
);
/*
    typedef logic[31:0][127:0] array_t ; 
    typedef logic[31:0][63:0] array_r ; 

    array_t rram_e = 'z ; 
    array_t rram_o = 'z ;

    array_r rd_en_e = '0 ;
    array_r rd_en_o = '0 ;

    logic [5:0] col ;
    logic [4:0] row ;
*/

endmodule