package comparator_pkg;
    typedef enum logic[7:0] {min, max, inf, inf_or_eq, eq, sup_or_eq, sup, neq} comparator_intr_e;
endpackage